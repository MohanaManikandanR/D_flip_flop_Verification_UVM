interface dff_interface();
  logic clk;
  logic rst;
  logic din;
  logic dout;
endinterface

  
